library verilog;
use verilog.vl_types.all;
entity decode_vlg_vec_tst is
end decode_vlg_vec_tst;
