library verilog;
use verilog.vl_types.all;
entity ersi_vlg_vec_tst is
end ersi_vlg_vec_tst;
